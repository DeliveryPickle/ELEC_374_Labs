library verilog;
use verilog.vl_types.all;
entity BusMux is
    port(
        R0Out           : in     vl_logic;
        R1Out           : in     vl_logic;
        R2Out           : in     vl_logic;
        R3Out           : in     vl_logic;
        R4Out           : in     vl_logic;
        R5Out           : in     vl_logic;
        R6Out           : in     vl_logic;
        R7Out           : in     vl_logic;
        R8Out           : in     vl_logic;
        R9Out           : in     vl_logic;
        R10Out          : in     vl_logic;
        R11Out          : in     vl_logic;
        R12Out          : in     vl_logic;
        R13Out          : in     vl_logic;
        R14Out          : in     vl_logic;
        R15Out          : in     vl_logic;
        hiOut           : in     vl_logic;
        loOut           : in     vl_logic;
        ZhiOut          : in     vl_logic;
        ZloOut          : in     vl_logic;
        PCout           : in     vl_logic;
        MDRout          : in     vl_logic;
        inPortout       : in     vl_logic;
        Cout            : in     vl_logic;
        busin0          : in     vl_logic_vector(31 downto 0);
        busin1          : in     vl_logic_vector(31 downto 0);
        busin2          : in     vl_logic_vector(31 downto 0);
        busin3          : in     vl_logic_vector(31 downto 0);
        busin4          : in     vl_logic_vector(31 downto 0);
        busin5          : in     vl_logic_vector(31 downto 0);
        busin6          : in     vl_logic_vector(31 downto 0);
        busin7          : in     vl_logic_vector(31 downto 0);
        busin8          : in     vl_logic_vector(31 downto 0);
        busin9          : in     vl_logic_vector(31 downto 0);
        busin10         : in     vl_logic_vector(31 downto 0);
        busin11         : in     vl_logic_vector(31 downto 0);
        busin12         : in     vl_logic_vector(31 downto 0);
        busin13         : in     vl_logic_vector(31 downto 0);
        busin14         : in     vl_logic_vector(31 downto 0);
        busin15         : in     vl_logic_vector(31 downto 0);
        businhi         : in     vl_logic_vector(31 downto 0);
        businlo         : in     vl_logic_vector(31 downto 0);
        businZhi        : in     vl_logic_vector(31 downto 0);
        businZlo        : in     vl_logic_vector(31 downto 0);
        businPC         : in     vl_logic_vector(31 downto 0);
        businMDR        : in     vl_logic_vector(31 downto 0);
        businInport     : in     vl_logic_vector(31 downto 0);
        csignextended   : in     vl_logic_vector(31 downto 0);
        busOut          : out    vl_logic_vector(31 downto 0)
    );
end BusMux;
