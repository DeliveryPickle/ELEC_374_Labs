library verilog;
use verilog.vl_types.all;
entity bus_tb is
end bus_tb;
